library verilog;
use verilog.vl_types.all;
entity LCD_Display_Controller_vlg_vec_tst is
end LCD_Display_Controller_vlg_vec_tst;
